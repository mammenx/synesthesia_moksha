parameter ACORTEX_I2C_BLK_CODE      = 0;
parameter ACORTEX_DRVR_BLK_CODE     = 1;
parameter ACORTEX_PCM_BFFR_CLK_CODE = 2;
