/*
 --------------------------------------------------------------------------
   Synesthesia-Moksha - Copyright (C) 2012 Gregory Matthew James.

   This file is part of Synesthesia-Moksha.

   Synesthesia-Moksha is free; you can redistribute it and/or modify
   it under the terms of the GNU General Public License as published by
   the Free Software Foundation; either version 3 of the License, or
   (at your option) any later version.

   Synesthesia-Moksha is distributed in the hope that it will be useful,
   but WITHOUT ANY WARRANTY; without even the implied warranty of
   MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE. See the
   GNU General Public License for more details.

   You should have received a copy of the GNU General Public License
   along with this program. If not, see <http://www.gnu.org/licenses/>.
 --------------------------------------------------------------------------
*/

/*
 --------------------------------------------------------------------------
 -- Project Code      : synesthesia_moksha
 -- Package Name      : syn_dsp_pkg
 -- Author            : mammenx
 -- Description       : This package contains DPI functions related to DSP
                        transforms.
 --------------------------------------------------------------------------
*/

package syn_dsp_pkg;

  import  syn_math_pkg::*;

  //import dpi task      C Name = SV function name
  import "DPI-C" pure function void syn_calc_fft(input int num_samples,input real data_in_arry[], inout real data_out_re_arry[], inout real data_out_im_arry[]);


endpackage : syn_dsp_pkg


/*
 --------------------------------------------------------------------------

 -- <Header>
 

 -- <Log>

[06-12-2014  05:46:09 PM][mammenx] Initial Commit

 --------------------------------------------------------------------------
*/


