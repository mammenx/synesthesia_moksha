// limbus.v

// Generated using ACDS version 13.1 162 at 2014.11.12.15:45:59

`timescale 1 ps / 1 ps
module limbus (
		input  wire        clk_clk,                                        //          clk.clk
		input  wire        reset_reset_n,                                  //        reset.reset_n
		output wire [0:0]  sram_bridge_sram_cntrlr_tcm_chipselect_n_out,   //  sram_bridge.sram_cntrlr_tcm_chipselect_n_out
		output wire [1:0]  sram_bridge_sram_cntrlr_tcm_byteenable_n_out,   //             .sram_cntrlr_tcm_byteenable_n_out
		output wire [18:0] sram_bridge_sram_cntrlr_tcm_address_out,        //             .sram_cntrlr_tcm_address_out
		output wire [0:0]  sram_bridge_sram_cntrlr_tcm_write_n_out,        //             .sram_cntrlr_tcm_write_n_out
		inout  wire [15:0] sram_bridge_sram_cntrlr_tcm_data_out,           //             .sram_cntrlr_tcm_data_out
		output wire [0:0]  sram_bridge_sram_cntrlr_tcm_outputenable_n_out, //             .sram_cntrlr_tcm_outputenable_n_out
		input  wire        uart_0_rxd,                                     //       uart_0.rxd
		output wire        uart_0_txd,                                     //             .txd
		output wire [17:0] cortex_s_address,                               //     cortex_s.address
		output wire        cortex_s_read,                                  //             .read
		input  wire [31:0] cortex_s_readdata,                              //             .readdata
		output wire        cortex_s_write,                                 //             .write
		output wire [31:0] cortex_s_writedata,                             //             .writedata
		input  wire        cortex_s_readdatavalid,                         //             .readdatavalid
		output wire        cortex_reset_reset,                             // cortex_reset.reset
		input  wire        cortex_irq_irq                                  //   cortex_irq.irq
	);

	wire         sram_cntrlr_tcm_chipselect_n_out;                           // sram_cntrlr:tcm_chipselect_n_out -> sram_pin_sharer:tcs0_chipselect_n_out
	wire         sram_cntrlr_tcm_grant;                                      // sram_pin_sharer:tcs0_grant -> sram_cntrlr:tcm_grant
	wire         sram_cntrlr_tcm_data_outen;                                 // sram_cntrlr:tcm_data_outen -> sram_pin_sharer:tcs0_data_outen
	wire         sram_cntrlr_tcm_outputenable_n_out;                         // sram_cntrlr:tcm_outputenable_n_out -> sram_pin_sharer:tcs0_outputenable_n_out
	wire         sram_cntrlr_tcm_request;                                    // sram_cntrlr:tcm_request -> sram_pin_sharer:tcs0_request
	wire  [15:0] sram_cntrlr_tcm_data_out;                                   // sram_cntrlr:tcm_data_out -> sram_pin_sharer:tcs0_data_out
	wire         sram_cntrlr_tcm_write_n_out;                                // sram_cntrlr:tcm_write_n_out -> sram_pin_sharer:tcs0_write_n_out
	wire  [18:0] sram_cntrlr_tcm_address_out;                                // sram_cntrlr:tcm_address_out -> sram_pin_sharer:tcs0_address_out
	wire  [15:0] sram_cntrlr_tcm_data_in;                                    // sram_pin_sharer:tcs0_data_in -> sram_cntrlr:tcm_data_in
	wire   [1:0] sram_cntrlr_tcm_byteenable_n_out;                           // sram_cntrlr:tcm_byteenable_n_out -> sram_pin_sharer:tcs0_byteenable_n_out
	wire   [0:0] sram_pin_sharer_tcm_sram_cntrlr_tcm_write_n_out_out;        // sram_pin_sharer:sram_cntrlr_tcm_write_n_out -> sram_bridge:tcs_sram_cntrlr_tcm_write_n_out
	wire  [15:0] sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_in;            // sram_bridge:tcs_sram_cntrlr_tcm_data_in -> sram_pin_sharer:sram_cntrlr_tcm_data_in
	wire   [0:0] sram_pin_sharer_tcm_sram_cntrlr_tcm_outputenable_n_out_out; // sram_pin_sharer:sram_cntrlr_tcm_outputenable_n_out -> sram_bridge:tcs_sram_cntrlr_tcm_outputenable_n_out
	wire         sram_pin_sharer_tcm_grant;                                  // sram_bridge:grant -> sram_pin_sharer:grant
	wire         sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_outen;         // sram_pin_sharer:sram_cntrlr_tcm_data_outen -> sram_bridge:tcs_sram_cntrlr_tcm_data_outen
	wire  [15:0] sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_out;           // sram_pin_sharer:sram_cntrlr_tcm_data_out -> sram_bridge:tcs_sram_cntrlr_tcm_data_out
	wire   [0:0] sram_pin_sharer_tcm_sram_cntrlr_tcm_chipselect_n_out_out;   // sram_pin_sharer:sram_cntrlr_tcm_chipselect_n_out -> sram_bridge:tcs_sram_cntrlr_tcm_chipselect_n_out
	wire         sram_pin_sharer_tcm_request;                                // sram_pin_sharer:request -> sram_bridge:request
	wire  [18:0] sram_pin_sharer_tcm_sram_cntrlr_tcm_address_out_out;        // sram_pin_sharer:sram_cntrlr_tcm_address_out -> sram_bridge:tcs_sram_cntrlr_tcm_address_out
	wire   [1:0] sram_pin_sharer_tcm_sram_cntrlr_tcm_byteenable_n_out_out;   // sram_pin_sharer:sram_cntrlr_tcm_byteenable_n_out -> sram_bridge:tcs_sram_cntrlr_tcm_byteenable_n_out
	wire         mm_interconnect_0_sram_cntrlr_uas_waitrequest;              // sram_cntrlr:uas_waitrequest -> mm_interconnect_0:sram_cntrlr_uas_waitrequest
	wire   [1:0] mm_interconnect_0_sram_cntrlr_uas_burstcount;               // mm_interconnect_0:sram_cntrlr_uas_burstcount -> sram_cntrlr:uas_burstcount
	wire  [15:0] mm_interconnect_0_sram_cntrlr_uas_writedata;                // mm_interconnect_0:sram_cntrlr_uas_writedata -> sram_cntrlr:uas_writedata
	wire  [18:0] mm_interconnect_0_sram_cntrlr_uas_address;                  // mm_interconnect_0:sram_cntrlr_uas_address -> sram_cntrlr:uas_address
	wire         mm_interconnect_0_sram_cntrlr_uas_lock;                     // mm_interconnect_0:sram_cntrlr_uas_lock -> sram_cntrlr:uas_lock
	wire         mm_interconnect_0_sram_cntrlr_uas_write;                    // mm_interconnect_0:sram_cntrlr_uas_write -> sram_cntrlr:uas_write
	wire         mm_interconnect_0_sram_cntrlr_uas_read;                     // mm_interconnect_0:sram_cntrlr_uas_read -> sram_cntrlr:uas_read
	wire  [15:0] mm_interconnect_0_sram_cntrlr_uas_readdata;                 // sram_cntrlr:uas_readdata -> mm_interconnect_0:sram_cntrlr_uas_readdata
	wire         mm_interconnect_0_sram_cntrlr_uas_debugaccess;              // mm_interconnect_0:sram_cntrlr_uas_debugaccess -> sram_cntrlr:uas_debugaccess
	wire         mm_interconnect_0_sram_cntrlr_uas_readdatavalid;            // sram_cntrlr:uas_readdatavalid -> mm_interconnect_0:sram_cntrlr_uas_readdatavalid
	wire   [1:0] mm_interconnect_0_sram_cntrlr_uas_byteenable;               // mm_interconnect_0:sram_cntrlr_uas_byteenable -> sram_cntrlr:uas_byteenable
	wire         cpu_instruction_master_waitrequest;                         // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [21:0] cpu_instruction_master_address;                             // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                            // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_data_master_waitrequest;                                // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                  // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [21:0] cpu_data_master_address;                                    // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire         cpu_data_master_write;                                      // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire         cpu_data_master_read;                                       // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                   // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_debugaccess;                                // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                 // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire  [15:0] mm_interconnect_0_uart_0_s1_writedata;                      // mm_interconnect_0:uart_0_s1_writedata -> uart_0:writedata
	wire   [2:0] mm_interconnect_0_uart_0_s1_address;                        // mm_interconnect_0:uart_0_s1_address -> uart_0:address
	wire         mm_interconnect_0_uart_0_s1_chipselect;                     // mm_interconnect_0:uart_0_s1_chipselect -> uart_0:chipselect
	wire         mm_interconnect_0_uart_0_s1_write;                          // mm_interconnect_0:uart_0_s1_write -> uart_0:write_n
	wire         mm_interconnect_0_uart_0_s1_read;                           // mm_interconnect_0:uart_0_s1_read -> uart_0:read_n
	wire  [15:0] mm_interconnect_0_uart_0_s1_readdata;                       // uart_0:readdata -> mm_interconnect_0:uart_0_s1_readdata
	wire         mm_interconnect_0_uart_0_s1_begintransfer;                  // mm_interconnect_0:uart_0_s1_begintransfer -> uart_0:begintransfer
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                     // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                       // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_chipselect;                    // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire         mm_interconnect_0_timer_0_s1_write;                         // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                      // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;              // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;             // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;  // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;     // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;        // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;          // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;            // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;              // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;               // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;           // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;        // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;         // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         irq_mapper_receiver0_irq;                                   // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                   // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                   // uart_0:irq -> irq_mapper:receiver2_irq
	wire  [31:0] cpu_d_irq_irq;                                              // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset_req;                         // rst_controller:reset_req -> [cpu:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                          // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	limbus_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~cortex_reset_reset),                                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	limbus_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~cortex_reset_reset),                                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	limbus_sram_cntrlr #(
		.TCM_ADDRESS_W                  (19),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (10),
		.TCM_WRITE_WAIT                 (10),
		.TCM_SETUP_WAIT                 (10),
		.TCM_DATA_HOLD                  (10),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) sram_cntrlr (
		.clk_clk                (clk_clk),                                         //   clk.clk
		.reset_reset            (cortex_reset_reset),                              // reset.reset
		.uas_address            (mm_interconnect_0_sram_cntrlr_uas_address),       //   uas.address
		.uas_burstcount         (mm_interconnect_0_sram_cntrlr_uas_burstcount),    //      .burstcount
		.uas_read               (mm_interconnect_0_sram_cntrlr_uas_read),          //      .read
		.uas_write              (mm_interconnect_0_sram_cntrlr_uas_write),         //      .write
		.uas_waitrequest        (mm_interconnect_0_sram_cntrlr_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid      (mm_interconnect_0_sram_cntrlr_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable         (mm_interconnect_0_sram_cntrlr_uas_byteenable),    //      .byteenable
		.uas_readdata           (mm_interconnect_0_sram_cntrlr_uas_readdata),      //      .readdata
		.uas_writedata          (mm_interconnect_0_sram_cntrlr_uas_writedata),     //      .writedata
		.uas_lock               (mm_interconnect_0_sram_cntrlr_uas_lock),          //      .lock
		.uas_debugaccess        (mm_interconnect_0_sram_cntrlr_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out        (sram_cntrlr_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_chipselect_n_out   (sram_cntrlr_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out (sram_cntrlr_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_request            (sram_cntrlr_tcm_request),                         //      .request
		.tcm_grant              (sram_cntrlr_tcm_grant),                           //      .grant
		.tcm_address_out        (sram_cntrlr_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out   (sram_cntrlr_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out           (sram_cntrlr_tcm_data_out),                        //      .data_out
		.tcm_data_outen         (sram_cntrlr_tcm_data_outen),                      //      .data_outen
		.tcm_data_in            (sram_cntrlr_tcm_data_in)                          //      .data_in
	);

	limbus_sram_pin_sharer sram_pin_sharer (
		.clk_clk                            (clk_clk),                                                    //   clk.clk
		.reset_reset                        (cortex_reset_reset),                                         // reset.reset
		.request                            (sram_pin_sharer_tcm_request),                                //   tcm.request
		.grant                              (sram_pin_sharer_tcm_grant),                                  //      .grant
		.sram_cntrlr_tcm_address_out        (sram_pin_sharer_tcm_sram_cntrlr_tcm_address_out_out),        //      .sram_cntrlr_tcm_address_out_out
		.sram_cntrlr_tcm_outputenable_n_out (sram_pin_sharer_tcm_sram_cntrlr_tcm_outputenable_n_out_out), //      .sram_cntrlr_tcm_outputenable_n_out_out
		.sram_cntrlr_tcm_byteenable_n_out   (sram_pin_sharer_tcm_sram_cntrlr_tcm_byteenable_n_out_out),   //      .sram_cntrlr_tcm_byteenable_n_out_out
		.sram_cntrlr_tcm_write_n_out        (sram_pin_sharer_tcm_sram_cntrlr_tcm_write_n_out_out),        //      .sram_cntrlr_tcm_write_n_out_out
		.sram_cntrlr_tcm_data_out           (sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_out),           //      .sram_cntrlr_tcm_data_out_out
		.sram_cntrlr_tcm_data_in            (sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_in),            //      .sram_cntrlr_tcm_data_out_in
		.sram_cntrlr_tcm_data_outen         (sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_outen),         //      .sram_cntrlr_tcm_data_out_outen
		.sram_cntrlr_tcm_chipselect_n_out   (sram_pin_sharer_tcm_sram_cntrlr_tcm_chipselect_n_out_out),   //      .sram_cntrlr_tcm_chipselect_n_out_out
		.tcs0_request                       (sram_cntrlr_tcm_request),                                    //  tcs0.request
		.tcs0_grant                         (sram_cntrlr_tcm_grant),                                      //      .grant
		.tcs0_address_out                   (sram_cntrlr_tcm_address_out),                                //      .address_out
		.tcs0_outputenable_n_out            (sram_cntrlr_tcm_outputenable_n_out),                         //      .outputenable_n_out
		.tcs0_byteenable_n_out              (sram_cntrlr_tcm_byteenable_n_out),                           //      .byteenable_n_out
		.tcs0_write_n_out                   (sram_cntrlr_tcm_write_n_out),                                //      .write_n_out
		.tcs0_data_out                      (sram_cntrlr_tcm_data_out),                                   //      .data_out
		.tcs0_data_in                       (sram_cntrlr_tcm_data_in),                                    //      .data_in
		.tcs0_data_outen                    (sram_cntrlr_tcm_data_outen),                                 //      .data_outen
		.tcs0_chipselect_n_out              (sram_cntrlr_tcm_chipselect_n_out)                            //      .chipselect_n_out
	);

	limbus_sram_bridge sram_bridge (
		.clk                                    (clk_clk),                                                    //   clk.clk
		.reset                                  (cortex_reset_reset),                                         // reset.reset
		.request                                (sram_pin_sharer_tcm_request),                                //   tcs.request
		.grant                                  (sram_pin_sharer_tcm_grant),                                  //      .grant
		.tcs_sram_cntrlr_tcm_chipselect_n_out   (sram_pin_sharer_tcm_sram_cntrlr_tcm_chipselect_n_out_out),   //      .sram_cntrlr_tcm_chipselect_n_out_out
		.tcs_sram_cntrlr_tcm_byteenable_n_out   (sram_pin_sharer_tcm_sram_cntrlr_tcm_byteenable_n_out_out),   //      .sram_cntrlr_tcm_byteenable_n_out_out
		.tcs_sram_cntrlr_tcm_address_out        (sram_pin_sharer_tcm_sram_cntrlr_tcm_address_out_out),        //      .sram_cntrlr_tcm_address_out_out
		.tcs_sram_cntrlr_tcm_write_n_out        (sram_pin_sharer_tcm_sram_cntrlr_tcm_write_n_out_out),        //      .sram_cntrlr_tcm_write_n_out_out
		.tcs_sram_cntrlr_tcm_data_out           (sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_out),           //      .sram_cntrlr_tcm_data_out_out
		.tcs_sram_cntrlr_tcm_data_outen         (sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_outen),         //      .sram_cntrlr_tcm_data_out_outen
		.tcs_sram_cntrlr_tcm_data_in            (sram_pin_sharer_tcm_sram_cntrlr_tcm_data_out_in),            //      .sram_cntrlr_tcm_data_out_in
		.tcs_sram_cntrlr_tcm_outputenable_n_out (sram_pin_sharer_tcm_sram_cntrlr_tcm_outputenable_n_out_out), //      .sram_cntrlr_tcm_outputenable_n_out_out
		.sram_cntrlr_tcm_chipselect_n_out       (sram_bridge_sram_cntrlr_tcm_chipselect_n_out),               //   out.sram_cntrlr_tcm_chipselect_n_out
		.sram_cntrlr_tcm_byteenable_n_out       (sram_bridge_sram_cntrlr_tcm_byteenable_n_out),               //      .sram_cntrlr_tcm_byteenable_n_out
		.sram_cntrlr_tcm_address_out            (sram_bridge_sram_cntrlr_tcm_address_out),                    //      .sram_cntrlr_tcm_address_out
		.sram_cntrlr_tcm_write_n_out            (sram_bridge_sram_cntrlr_tcm_write_n_out),                    //      .sram_cntrlr_tcm_write_n_out
		.sram_cntrlr_tcm_data_out               (sram_bridge_sram_cntrlr_tcm_data_out),                       //      .sram_cntrlr_tcm_data_out
		.sram_cntrlr_tcm_outputenable_n_out     (sram_bridge_sram_cntrlr_tcm_outputenable_n_out)              //      .sram_cntrlr_tcm_outputenable_n_out
	);

	limbus_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~cortex_reset_reset),                     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	limbus_uart_0 uart_0 (
		.clk           (clk_clk),                                   //                 clk.clk
		.reset_n       (~cortex_reset_reset),                       //               reset.reset_n
		.address       (mm_interconnect_0_uart_0_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_0_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_0_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_0_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_0_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_0_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_0_s1_readdata),      //                    .readdata
		.dataavailable (),                                          //                    .dataavailable
		.readyfordata  (),                                          //                    .readyfordata
		.rxd           (uart_0_rxd),                                // external_connection.export
		.txd           (uart_0_txd),                                //                    .export
		.irq           (irq_mapper_receiver2_irq)                   //                 irq.irq
	);

	limbus_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~cortex_reset_reset),                            //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	limbus_mm_interconnect_0 mm_interconnect_0 (
		.clk_100_clk_clk                         (clk_clk),                                                   //                       clk_100_clk.clk
		.cpu_reset_n_reset_bridge_in_reset_reset (cortex_reset_reset),                                        // cpu_reset_n_reset_bridge_in_reset.reset
		.cpu_data_master_address                 (cpu_data_master_address),                                   //                   cpu_data_master.address
		.cpu_data_master_waitrequest             (cpu_data_master_waitrequest),                               //                                  .waitrequest
		.cpu_data_master_byteenable              (cpu_data_master_byteenable),                                //                                  .byteenable
		.cpu_data_master_read                    (cpu_data_master_read),                                      //                                  .read
		.cpu_data_master_readdata                (cpu_data_master_readdata),                                  //                                  .readdata
		.cpu_data_master_write                   (cpu_data_master_write),                                     //                                  .write
		.cpu_data_master_writedata               (cpu_data_master_writedata),                                 //                                  .writedata
		.cpu_data_master_debugaccess             (cpu_data_master_debugaccess),                               //                                  .debugaccess
		.cpu_instruction_master_address          (cpu_instruction_master_address),                            //            cpu_instruction_master.address
		.cpu_instruction_master_waitrequest      (cpu_instruction_master_waitrequest),                        //                                  .waitrequest
		.cpu_instruction_master_read             (cpu_instruction_master_read),                               //                                  .read
		.cpu_instruction_master_readdata         (cpu_instruction_master_readdata),                           //                                  .readdata
		.cortex_s0_address                       (cortex_s_address),                                          //                         cortex_s0.address
		.cortex_s0_write                         (cortex_s_write),                                            //                                  .write
		.cortex_s0_read                          (cortex_s_read),                                             //                                  .read
		.cortex_s0_readdata                      (cortex_s_readdata),                                         //                                  .readdata
		.cortex_s0_writedata                     (cortex_s_writedata),                                        //                                  .writedata
		.cortex_s0_readdatavalid                 (cortex_s_readdatavalid),                                    //                                  .readdatavalid
		.cpu_jtag_debug_module_address           (mm_interconnect_0_cpu_jtag_debug_module_address),           //             cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write             (mm_interconnect_0_cpu_jtag_debug_module_write),             //                                  .write
		.cpu_jtag_debug_module_read              (mm_interconnect_0_cpu_jtag_debug_module_read),              //                                  .read
		.cpu_jtag_debug_module_readdata          (mm_interconnect_0_cpu_jtag_debug_module_readdata),          //                                  .readdata
		.cpu_jtag_debug_module_writedata         (mm_interconnect_0_cpu_jtag_debug_module_writedata),         //                                  .writedata
		.cpu_jtag_debug_module_byteenable        (mm_interconnect_0_cpu_jtag_debug_module_byteenable),        //                                  .byteenable
		.cpu_jtag_debug_module_waitrequest       (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),       //                                  .waitrequest
		.cpu_jtag_debug_module_debugaccess       (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),       //                                  .debugaccess
		.jtag_uart_avalon_jtag_slave_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //       jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                  .write
		.jtag_uart_avalon_jtag_slave_read        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                  .read
		.jtag_uart_avalon_jtag_slave_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                  .readdata
		.jtag_uart_avalon_jtag_slave_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                  .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.sram_cntrlr_uas_address                 (mm_interconnect_0_sram_cntrlr_uas_address),                 //                   sram_cntrlr_uas.address
		.sram_cntrlr_uas_write                   (mm_interconnect_0_sram_cntrlr_uas_write),                   //                                  .write
		.sram_cntrlr_uas_read                    (mm_interconnect_0_sram_cntrlr_uas_read),                    //                                  .read
		.sram_cntrlr_uas_readdata                (mm_interconnect_0_sram_cntrlr_uas_readdata),                //                                  .readdata
		.sram_cntrlr_uas_writedata               (mm_interconnect_0_sram_cntrlr_uas_writedata),               //                                  .writedata
		.sram_cntrlr_uas_burstcount              (mm_interconnect_0_sram_cntrlr_uas_burstcount),              //                                  .burstcount
		.sram_cntrlr_uas_byteenable              (mm_interconnect_0_sram_cntrlr_uas_byteenable),              //                                  .byteenable
		.sram_cntrlr_uas_readdatavalid           (mm_interconnect_0_sram_cntrlr_uas_readdatavalid),           //                                  .readdatavalid
		.sram_cntrlr_uas_waitrequest             (mm_interconnect_0_sram_cntrlr_uas_waitrequest),             //                                  .waitrequest
		.sram_cntrlr_uas_lock                    (mm_interconnect_0_sram_cntrlr_uas_lock),                    //                                  .lock
		.sram_cntrlr_uas_debugaccess             (mm_interconnect_0_sram_cntrlr_uas_debugaccess),             //                                  .debugaccess
		.sysid_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),             //               sysid_control_slave.address
		.sysid_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata),            //                                  .readdata
		.timer_0_s1_address                      (mm_interconnect_0_timer_0_s1_address),                      //                        timer_0_s1.address
		.timer_0_s1_write                        (mm_interconnect_0_timer_0_s1_write),                        //                                  .write
		.timer_0_s1_readdata                     (mm_interconnect_0_timer_0_s1_readdata),                     //                                  .readdata
		.timer_0_s1_writedata                    (mm_interconnect_0_timer_0_s1_writedata),                    //                                  .writedata
		.timer_0_s1_chipselect                   (mm_interconnect_0_timer_0_s1_chipselect),                   //                                  .chipselect
		.uart_0_s1_address                       (mm_interconnect_0_uart_0_s1_address),                       //                         uart_0_s1.address
		.uart_0_s1_write                         (mm_interconnect_0_uart_0_s1_write),                         //                                  .write
		.uart_0_s1_read                          (mm_interconnect_0_uart_0_s1_read),                          //                                  .read
		.uart_0_s1_readdata                      (mm_interconnect_0_uart_0_s1_readdata),                      //                                  .readdata
		.uart_0_s1_writedata                     (mm_interconnect_0_uart_0_s1_writedata),                     //                                  .writedata
		.uart_0_s1_begintransfer                 (mm_interconnect_0_uart_0_s1_begintransfer),                 //                                  .begintransfer
		.uart_0_s1_chipselect                    (mm_interconnect_0_uart_0_s1_chipselect)                     //                                  .chipselect
	);

	limbus_irq_mapper irq_mapper (
		.clk           (clk_clk),                  //       clk.clk
		.reset         (cortex_reset_reset),       // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.receiver3_irq (cortex_irq_irq),           // receiver3.irq
		.sender_irq    (cpu_d_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (cortex_reset_reset),                 // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
