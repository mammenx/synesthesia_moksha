parameter SYS_MEM_HST_ACC_STATUS_REG  = 0;
parameter SYS_MEM_HST_ACC_ADDR_REG    = 1;
parameter SYS_MEM_HST_ACC_DATA_REG    = 2;
