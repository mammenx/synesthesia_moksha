parameter RST_CNTRL_REG_ADDR = 0;
