//Block Code
parameter ACORTEX_BLK               = 0;
parameter FGYRUS_BLK                = 1;
parameter RST_SYNC_BLK              = 2;
parameter SYS_MEM_MNGR_BLK          = 3;
//parameter VCORTEX_BLK               = 1;
