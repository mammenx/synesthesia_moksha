parameter RST_CNTRL_REG_ADDR        = 0;
parameter RST_CNTRL_NUM_RESETS_ADDR = 1;
