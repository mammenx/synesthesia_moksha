parameter SYS_MEM_ARB_STATUS_REG    = 0;
