parameter ADV7513_CNTRLR_CONFIG_REG     = 0;
parameter ADV7513_CNTRLR_STATUS_REG     = 1;
parameter ADV7513_CNTRLR_LBFFR_OCC_REG  = 2;
