parameter I2C_ADDR_REG_ADDR         = 0;
parameter I2C_CLK_DIV_REG_ADDR      = 1;
parameter I2C_CONFIG_REG_ADDR       = 2;
parameter I2C_STATUS_REG_ADDR       = 3;
parameter I2C_FSM_REG_ADDR          = 4;
parameter I2C_DATA_CACHE_BASE_ADDR  = 5;
