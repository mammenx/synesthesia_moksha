//Block Code
parameter ACORTEX_BLK               = 0;
parameter RST_SYNC_BLK              = 1;
//parameter VCORTEX_BLK               = 1;
//parameter FGYRUS_BLK                = 2;
