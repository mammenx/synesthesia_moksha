parameter SYS_MEM_INTF_ARB_BLK_CODE   = 0;
parameter SYS_MEM_INTF_PART_BLK_CODE  = 1;
