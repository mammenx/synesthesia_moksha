parameter GRAPHEME_LB_BLK_CODE        = 0;
parameter GRAPHEME_HST_ACC_BLK_CODE   = 1;
