parameter SSM2603_DRVR_CONFIG_REG_ADDR    = 0;
parameter SSM2603_DRVR_STATUS_REG_ADDR    = 1;
parameter SSM2603_DRVR_BCLK_DIV_REG_ADDR  = 2;
parameter SSM2603_DRVR_FS_VAL_REG_ADDR    = 3;
